
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
USE ieee.numeric_std.ALL;


entity RF is
    port (
          RD : in std_logic_vector(5 downto 0);
          DWR   : in std_logic_vector(31 downto 0);
			 RS1   : in std_logic_vector(5 downto 0);
			 RS2   : in std_logic_vector(5 downto 0);
          CRS1   : out std_logic_vector(31 downto 0);
			 CRS2   : out std_logic_vector(31 downto 0);
			 CRD: out std_logic_vector(31 downto 0);
			 rst: in std_logic;
			 we: in std_logic
			 );
end RF;

architecture syn of RF is
    type ram_type is array (0 to 39) of std_logic_vector (31 downto 0);
    signal RAM: ram_type;
	 signal rdaux: std_logic_vector(5 downto 0);

begin
	 rdaux <= rd;
    process (RDaux,RS1,RS2,rst,we)
    begin
			RAM(0) <= "00000000000000000000000000000000";
			CRS1 <= RAM(to_integer(unsigned(RS1)));
			CRS2 <= RAM(to_integer(unsigned(RS2)));
			CRD <=  RAM(to_integer(unsigned(RD)));

			if(RD /= "000000" and we = '1') then
				RAM(conv_integer(RDaux)) <= DWR;
			end if;
        if rst = '1' then
				RAM(0) <= "00000000000000000000000000000000";
				RAM(1) <= "00000000000000000000000000000000";
				RAM(2) <= "00000000000000000000000000000000";
				RAM(3) <= "00000000000000000000000000000000";
				RAM(4) <= "00000000000000000000000000000000";
				RAM(5) <= "00000000000000000000000000000000";
				RAM(6) <= "00000000000000000000000000000000";
				RAM(7) <= "00000000000000000000000000000000";
				RAM(8) <= "00000000000000000000000000000000";
				RAM(9) <= "00000000000000000000000000000000";
				RAM(10) <= "00000000000000000000000000000000";
				RAM(11) <= "00000000000000000000000000000000";
				RAM(12) <= "00000000000000000000000000000000";
				RAM(13) <= "00000000000000000000000000000000";
				RAM(14) <= "00000000000000000000000000000000";
				RAM(15) <= "00000000000000000000000000000000";
				RAM(16) <= "00000000000000000000000000000000";
				RAM(17) <= "00000000000000000000000000000000";
				RAM(18) <= "00000000000000000000000000000000";
				RAM(19) <= "00000000000000000000000000000000";
				RAM(20) <= "00000000000000000000000000000000";
				RAM(21) <= "00000000000000000000000000000000";
				RAM(22) <= "00000000000000000000000000000000";
				RAM(23) <= "00000000000000000000000000000000";
				RAM(24) <= "00000000000000000000000000000000";
				RAM(25) <= "00000000000000000000000000000000";
				RAM(26) <= "00000000000000000000000000000000";
				RAM(27) <= "00000000000000000000000000000000";
				RAM(28) <= "00000000000000000000000000000000";
				RAM(29) <= "00000000000000000000000000000000";
				RAM(30) <= "00000000000000000000000000000000";
				RAM(31) <= "00000000000000000000000000000000";
				RAM(32) <= "00000000000000000000000000000000";	
				RAM(33) <= "00000000000000000000000000000000";	
				RAM(34) <= "00000000000000000000000000000000";	
				RAM(35) <= "00000000000000000000000000000000";	
				RAM(36) <= "00000000000000000000000000000000";	
				RAM(37) <= "00000000000000000000000000000000";	
				RAM(38) <= "00000000000000000000000000000000";	
				RAM(39) <= "00000000000000000000000000000000";	
        end if;
    end process;

end syn;