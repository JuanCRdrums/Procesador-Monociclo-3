library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity instructionMemory is
port (rst : in  STD_LOGIC;
      EN : in std_logic;
      ADDR : in std_logic_vector(31 downto 0);
      DATA : out std_logic_vector(31 downto 0));
end instructionMemory;

architecture syn of instructionMemory is
    type rom_type is array (0 to 63) of std_logic_vector (31 downto 0);                 
    signal ROM : rom_type:= ("10100000000100000010000000000101", "10100100000100000010000000000000","10000001110000000010000000000101", "10100010000100000010000000001000", "00000001000000000000000000000000", "10000000101000001100000000010001",
                             "00000010100000000000000000000101", "00000001000000000000000000000000","10000110000000000111000000000001", "01111111111111111111111111111100", "10100000000001000000000000010000", "10010000000100000000000000010000",
                             "00000001000000000000000000000000", "00000001000000000000000000000000","00000001000000000000000000000000", "00000001000000000000000000000000", "00000001000000000000000000000000", "00000001000000000000000000000000",
                             "00000001000000000000000000000000", "00000001000000000000000000000000","00000001000000000000000000000000", "00000001000000000000000000000000", "00000001000000000000000000000000", "00000001000000000000000000000000",
                             "00000001000000000000000000000000", "00000001000000000000000000000000","00000001000000000000000000000000", "00000001000000000000000000000000", "00000001000000000000000000000000", "00000001000000000000000000000000",
                             "00000001000000000000000000000000", "00000001000000000000000000000000","00000001000000000000000000000000", "00000001000000000000000000000000", "00000001000000000000000000000000", "00000001000000000000000000000000",
                             "00000001000000000000000000000000", "00000001000000000000000000000000","00000001000000000000000000000000", "00000001000000000000000000000000", "00000001000000000000000000000000", "00000001000000000000000000000000",
                             "00000001000000000000000000000000", "00000001000000000000000000000000","00000001000000000000000000000000", "00000001000000000000000000000000", "00000001000000000000000000000000", "00000001000000000000000000000000",
                             "00000001000000000000000000000000", "00000001000000000000000000000000","00000001000000000000000000000000", "00000001000000000000000000000000", "00000001000000000000000000000000", "00000001000000000000000000000000",
                             "00000001000000000000000000000000", "00000001000000000000000000000000","00000001000000000000000000000000", "00000001000000000000000000000000", "00000001000000000000000000000000", "00000001000000000000000000000000",
                             "00000001000000000000000000000000", "00000001000000000000000000000000","00000001000000000000000000000000", "00000001000000000000000000000000" );                        



begin


	 
	
process(rst,ADDR)
	begin
	
	if rst = '1' then
		DATA<="00000000000000000000000000000000";
	else
		DATA <= ROM(conv_integer(ADDR(5 downto 0))); 
	end if;

end process;

end syn;